library verilog;
use verilog.vl_types.all;
entity SYNC_signal_vlg_vec_tst is
end SYNC_signal_vlg_vec_tst;
