-- HACER MAQUINA DE ESTADOS