library verilog;
use verilog.vl_types.all;
entity mainVGA_vlg_vec_tst is
end mainVGA_vlg_vec_tst;
